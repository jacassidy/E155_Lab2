// James Kaden Cassidy kacassidy@hmc.edu 9/7/2025
